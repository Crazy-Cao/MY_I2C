
`define SYS_CLK_100M
//`define	SYS_CLK_50M