
`define SYS_CLK_100M
//`define	SYS_CLK_50M
`define I2C_SPEED_CLK_100K
//`define IWC_SPEED_CLK_400K
